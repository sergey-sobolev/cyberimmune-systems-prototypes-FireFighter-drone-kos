component ffd.MovementActions

endpoints {
    actions: ffd.MovementActions
}
