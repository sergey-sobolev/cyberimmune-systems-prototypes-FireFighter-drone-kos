component ffd.CCUActions

endpoints {
    actions: ffd.CCUActions
}
