component ffd.CommunicationOutside

endpoints {
    startedat: ffd.CommunicationOutside
}
