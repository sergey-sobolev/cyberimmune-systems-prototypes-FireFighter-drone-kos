component ffd.CCUActions

endpoints {
    coordinates: ffd.CCUActions
}
