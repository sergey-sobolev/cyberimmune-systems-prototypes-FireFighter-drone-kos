component ffd.SituationActions

endpoints {
    actions: ffd.SituationActions
}
