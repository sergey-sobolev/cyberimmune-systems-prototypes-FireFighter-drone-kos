component ffd.AggregationCoordinates

endpoints {
    coordinates: ffd.AggregationCoordinates
}
