component ffd.ExtinguishingActions

endpoints {
    actions: ffd.ExtinguishingActions
}
