component ffd.FMACActions

endpoints {
    actions: ffd.FMACActions
}
