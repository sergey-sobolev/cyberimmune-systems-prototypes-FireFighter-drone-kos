component ffd.NavigationCoordinates

endpoints {
    coordinates: ffd.NavigationCoordinates
}
