component ffd.EAICActions

endpoints {
    actions: ffd.EAICActions
}
